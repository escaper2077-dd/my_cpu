module(

);

endmodule
